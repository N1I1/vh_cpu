`define ALU_ADD     4'b0000
`define ALU_SUB     4'b0001
`define ALU_AND     4'b0010
`define ALU_OR      4'b0011
`define ALU_XOR     4'b0100
`define ALU_SLL     4'b0101 // Shift left logical
`define ALU_SRL     4'b0110 // Shift right logical
`define ALU_SRA     4'b0111 // Shift right arithmetic
`define ALU_SLT     4'b1000 // Set less than
`define ALU_SLTU    4'b1001 // Set less than unsigned
`define ALU_COPY1   4'b1010 // Copy input 1 to output
`define ALU_COPY2   4'b1011 // Copy input 2 to output
`define ALU_MUL     4'b1100 // Multiply
`define ALU_JALR    4'b1101 // Jump and link register
`define ALU_CSRRC   4'b1110
`define ALU_XXX     4'bzzzz 