`include "../include/common.vh"

module pipe_mem_wb_reg(
    input clk,
    input rst,
    input mem_wb_en,
    input mem_wb_stall,
    input ...
    output reg ...
    );
    always @(posedge clk) begin
        if (rst) begin
            
        end else if (mem_wb_en) begin
            
        end else begin
            
        end
    end
endmodule