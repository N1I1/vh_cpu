`include "opcode.vh"
`include "alu.vh"
`include "../Color.vh"

`define ARCH_WIDTH 64
`define ALU_OP_WIDTH 4
`define ARCH "riscv64"
