`include "../include/common.vh"

module pipe_id_ex_reg(
    input clk,
    input rst,
    input id_ex_en,
    input id_ex_stall,
    input ...
    output reg ...
    );
    always @(posedge clk) begin
        if (rst) begin
            
        end else if (id_ex_en) begin
            
        end else begin
            
        end
    end
endmodule