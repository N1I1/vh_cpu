`include "opcode.vh"
`include "alu.vh"
`include "../Color.vh"
`include "func.vh"

`define ARCH_WIDTH 64
`define ALU_OP_WIDTH 4
`define ARCH "riscv64"

`define INSTR_WIDTH 32
`define INSTR_MEM_SIZE 65535
`define INSTR_MEM_WIDTH 64

`define DATA_WIDTH 64
`define DATA_MEM_SIZE 8192
`define DATA_MEM_WIDTH 64

`define DATA_WIDTH_8 3'd0
`define DATA_WIDTH_16 3'd1
`define DATA_WIDTH_32 3'd2
`define DATA_WIDTH_64 3'd3