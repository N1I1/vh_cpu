`include "../include/common.vh"

module mux8_1(
    input   wire    [2:0]   sel,
    input   wire    [`ARCH_WIDTH-1:0]  a,
    input   wire    [`ARCH_WIDTH-1:0]  b,
    input   wire    [`ARCH_WIDTH-1:0]  c,
    input   wire    [`ARCH_WIDTH-1:0]  d,
    input   wire    [`ARCH_WIDTH-1:0]  e,
    input   wire    [`ARCH_WIDTH-1:0]  f,
    input   wire    [`ARCH_WIDTH-1:0]  g,
    input   wire    [`ARCH_WIDTH-1:0]  h,
    output  reg     [`ARCH_WIDTH-1:0]  out
);

    always @(*) begin
        case(sel)
            3'b000: out = a;
            3'b001: out = b;
            3'b010: out = c;
            3'b011: out = d;
            3'b100: out = e;
            3'b101: out = f;
            3'b110: out = g;
            3'b111: out = h;
        endcase
    end

endmodule