`define ARCH_WIDTH 32
`define ALU_OP_WIDTH 5
`define ARCH "riscv32"