`include "../include/common.vh"

module pipe_ex_mem_reg(
    input clk,
    input rst,
    input ex_mem_en,
    input ex_mem_stall,
    input ...
    output reg ...
    );
    always @(posedge clk) begin
        if (rst) begin
            
        end else if (ex_mem_en) begin
            
        end else begin
            
        end
    end
endmodule